library verilog;
use verilog.vl_types.all;
entity ShiftLight_vlg_vec_tst is
end ShiftLight_vlg_vec_tst;
